*** SPICE deck for cell INVERTER{lay} from library MOSIS_SUBM_PADS_C5
*** Created on Sal Ara 12, 2023 13:55:25
*** Last revised on Sal Ara 12, 2023 15:00:23
*** Written on Sal Ara 12, 2023 15:00:28 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:\Users\mehme\OneDrive\tsmc018.txt

*** TOP LEVEL CELL: INVERTER{lay}
Mnmos@0 gnd a out gnd N L=0.6U W=0.9U AS=2.52P AD=2.52P PS=6.6U PD=6.6U
Mpmos@0 out a vdd vdd P L=0.6U W=0.9U AS=2.52P AD=2.52P PS=6.6U PD=6.6U

* Spice Code nodes in cell cell 'INVERTER{lay}'
vdd vdd 0 DC 5
va a 0 DC 0
vgnd gnd 0 DC 0
.dc va 5 5 5
.END
