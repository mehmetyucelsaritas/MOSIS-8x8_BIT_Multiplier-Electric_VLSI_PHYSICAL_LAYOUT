*** SPICE deck for cell HALF_ADDER{lay} from library MOSIS_SUBM_PADS_C5
*** Created on Sal Ara 12, 2023 18:23:00
*** Last revised on Sal Ara 12, 2023 20:33:02
*** Written on Sal Ara 12, 2023 20:33:05 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:\Users\mehme\OneDrive\tsmc018.txt

*** SUBCIRCUIT MOSIS_SUBM_PADS_C5__INVERTER FROM CELL INVERTER{lay}
.SUBCKT MOSIS_SUBM_PADS_C5__INVERTER a gnd out vdd
Mnmos@0 gnd a out gnd N L=0.6U W=0.9U AS=5.265P AD=2.52P PS=13.2U PD=6.6U
Mpmos@0 out a vdd vdd P L=0.6U W=0.9U AS=2.52P AD=5.265P PS=6.6U PD=13.2U
.ENDS MOSIS_SUBM_PADS_C5__INVERTER

*** SUBCIRCUIT MOSIS_SUBM_PADS_C5__AND_GATE FROM CELL AND_GATE{lay}
.SUBCKT MOSIS_SUBM_PADS_C5__AND_GATE a b gnd out vdd
XINVERTER@1 net@2 gnd out vdd MOSIS_SUBM_PADS_C5__INVERTER
Mnmos@2 net@0 b gnd gnd N L=0.6U W=0.9U AS=4.77P AD=0.742P PS=12.6U PD=2.55U
Mnmos@3 net@2 a net@0 gnd N L=0.6U W=0.9U AS=0.742P AD=3.735P PS=2.55U PD=9.3U
Mpmos@0 vdd b net@2 vdd P L=0.6U W=0.9U AS=3.735P AD=1.395P PS=9.3U PD=3.6U
Mpmos@1 net@2 a vdd vdd P L=0.6U W=0.9U AS=1.395P AD=3.735P PS=3.6U PD=9.3U
.ENDS MOSIS_SUBM_PADS_C5__AND_GATE

*** SUBCIRCUIT MOSIS_SUBM_PADS_C5__XOR_GATE FROM CELL XOR_GATE{lay}
.SUBCKT MOSIS_SUBM_PADS_C5__XOR_GATE a b gnd out vdd
XINVERTER@0 b gnd net@39 vdd MOSIS_SUBM_PADS_C5__INVERTER
XINVERTER@1 a gnd net@42 vdd MOSIS_SUBM_PADS_C5__INVERTER
Mnmos@0 net@1 a gnd gnd N L=0.6U W=0.9U AS=3.847P AD=0.742P PS=10.05U PD=2.55U
Mnmos@1 out b net@1 gnd N L=0.6U W=0.9U AS=0.742P AD=1.395P PS=2.55U PD=3.6U
Mnmos@2 net@4 net@39 out gnd N L=0.6U W=0.9U AS=1.395P AD=0.742P PS=3.6U PD=2.55U
Mnmos@3 gnd net@42 net@4 gnd N L=0.6U W=0.9U AS=0.742P AD=3.847P PS=2.55U PD=10.05U
Mpmos@0 vdd a net@6 vdd P L=0.6U W=0.9U AS=2.768P AD=1.395P PS=6.9U PD=3.6U
Mpmos@1 net@6 b vdd vdd P L=0.6U W=0.9U AS=1.395P AD=2.768P PS=3.6U PD=6.9U
Mpmos@2 out net@39 net@6 vdd P L=0.6U W=0.9U AS=2.768P AD=1.395P PS=6.9U PD=3.6U
Mpmos@3 net@6 net@42 out vdd P L=0.6U W=0.9U AS=1.395P AD=2.768P PS=3.6U PD=6.9U
.ENDS MOSIS_SUBM_PADS_C5__XOR_GATE

*** TOP LEVEL CELL: HALF_ADDER{lay}
XAND_GATE@8 a b gnd CARRY vdd MOSIS_SUBM_PADS_C5__AND_GATE
XXOR_GATE@2 a b gnd SUM vdd MOSIS_SUBM_PADS_C5__XOR_GATE

* Spice Code nodes in cell cell 'HALF_ADDER{lay}'
vdd vdd 0 dc 5
va a 0 dc 5
vb b 0 dc 5
.dc va 5 5 5 vb 5 5 5 
.END
