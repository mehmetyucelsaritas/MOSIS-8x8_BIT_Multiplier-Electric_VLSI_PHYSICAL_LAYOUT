*** SPICE deck for cell OR_GATE{lay} from library MOSIS_SUBM_PADS_C5
*** Created on Sal Ara 12, 2023 15:31:31
*** Last revised on Sal Ara 12, 2023 20:16:15
*** Written on Sal Ara 12, 2023 20:16:18 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:\Users\mehme\OneDrive\tsmc018.txt

*** SUBCIRCUIT MOSIS_SUBM_PADS_C5__INVERTER FROM CELL INVERTER{lay}
.SUBCKT MOSIS_SUBM_PADS_C5__INVERTER a gnd out vdd
Mnmos@0 gnd a out gnd N L=0.6U W=0.9U AS=5.265P AD=2.52P PS=13.2U PD=6.6U
Mpmos@0 out a vdd vdd P L=0.6U W=0.9U AS=2.52P AD=5.265P PS=6.6U PD=13.2U
.ENDS MOSIS_SUBM_PADS_C5__INVERTER

*** TOP LEVEL CELL: OR_GATE{lay}
XINVERTER@0 net@2 gnd out vdd MOSIS_SUBM_PADS_C5__INVERTER
Mnmos@0 net@2 a gnd gnd N L=0.6U W=0.9U AS=1.395P AD=3.27P PS=3.6U PD=8.6U
Mnmos@1 gnd b net@2 gnd N L=0.6U W=0.9U AS=3.27P AD=1.395P PS=8.6U PD=3.6U
Mpmos@0 net@0 b vdd vdd P L=0.6U W=0.9U AS=5.76P AD=0.742P PS=13.8U PD=2.55U
Mpmos@1 net@2 a net@0 vdd P L=0.6U W=0.9U AS=0.742P AD=3.27P PS=2.55U PD=8.6U

* Spice Code nodes in cell cell 'OR_GATE{lay}'
vdd vdd 0 dc 5
va a 0 dc 5
vb b 0 dc 5
.dc vdd 5 5 5 va 0 0 5 vb 0 0 5 vgnd 0 0 0
.END
