*** SPICE deck for cell XOR_GATE_trans{lay} from library MOSIS_SUBM_PADS_C5
*** Created on Sal Ara 12, 2023 15:56:57
*** Last revised on Sal Ara 12, 2023 16:35:04
*** Written on Sal Ara 12, 2023 16:35:06 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:\Users\mehme\OneDrive\tsmc018.txt

*** SUBCIRCUIT MOSIS_SUBM_PADS_C5__INVERTER FROM CELL INVERTER{lay}
.SUBCKT MOSIS_SUBM_PADS_C5__INVERTER a gnd out vdd
Mnmos@0 gnd a out gnd N L=0.6U W=0.9U AS=2.52P AD=2.52P PS=6.6U PD=6.6U
Mpmos@0 out a vdd vdd P L=0.6U W=0.9U AS=2.52P AD=2.52P PS=6.6U PD=6.6U
.ENDS MOSIS_SUBM_PADS_C5__INVERTER

*** TOP LEVEL CELL: XOR_GATE_trans{lay}
XINVERTER@0 a net@4 out b MOSIS_SUBM_PADS_C5__INVERTER
XINVERTER@2 b gnd net@4 vdd MOSIS_SUBM_PADS_C5__INVERTER
Mnmos@0 a net@4 out gnd N L=0.6U W=0.9U AS=2.52P AD=2.52P PS=6.6U PD=6.6U
Mpmos@0 a b out vdd P L=0.6U W=0.9U AS=2.52P AD=2.52P PS=6.6U PD=6.6U

* Spice Code nodes in cell cell 'XOR_GATE_trans{lay}'
vdd vdd 0 dc 5
vgnd gnd 0 dc 0
va a 0 dc 0
vb b 0 dc 0
.dc va 5 5 5 vb 0 0 5 vdd 5 5 5 vgnd 0 0 5
.END
